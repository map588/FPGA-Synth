library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

package midi_lut_pkg is
    type phase_inc_lut_type is array (0 to 127) of std_logic_vector(24 downto 0);
    constant midi_phase_inc_lut : phase_inc_lut_type;
end package midi_lut_pkg;

package body midi_lut_pkg is
    constant midi_phase_inc_lut: phase_inc_lut_type := (
        X"000594",  -- MIDI Note 0, Freq 8.18 Hz
        X"0005E9",  -- MIDI Note 1, Freq 8.66 Hz
        X"000643",  -- MIDI Note 2, Freq 9.18 Hz
        X"0006A3",  -- MIDI Note 3, Freq 9.72 Hz
        X"000708",  -- MIDI Note 4, Freq 10.30 Hz
        X"000773",  -- MIDI Note 5, Freq 10.91 Hz
        X"0007E4",  -- MIDI Note 6, Freq 11.56 Hz
        X"00085C",  -- MIDI Note 7, Freq 12.25 Hz
        X"0008DC",  -- MIDI Note 8, Freq 12.98 Hz
        X"000962",  -- MIDI Note 9, Freq 13.75 Hz
        X"0009F1",  -- MIDI Note 10, Freq 14.57 Hz
        X"000A89",  -- MIDI Note 11, Freq 15.43 Hz
        X"000B29",  -- MIDI Note 12, Freq 16.35 Hz
        X"000BD3",  -- MIDI Note 13, Freq 17.32 Hz
        X"000C87",  -- MIDI Note 14, Freq 18.35 Hz
        X"000D46",  -- MIDI Note 15, Freq 19.45 Hz
        X"000E10",  -- MIDI Note 16, Freq 20.60 Hz
        X"000EE6",  -- MIDI Note 17, Freq 21.83 Hz
        X"000FC9",  -- MIDI Note 18, Freq 23.12 Hz
        X"0010B9",  -- MIDI Note 19, Freq 24.50 Hz
        X"0011B8",  -- MIDI Note 20, Freq 25.96 Hz
        X"0012C5",  -- MIDI Note 21, Freq 27.50 Hz
        X"0013E3",  -- MIDI Note 22, Freq 29.14 Hz
        X"001512",  -- MIDI Note 23, Freq 30.87 Hz
        X"001653",  -- MIDI Note 24, Freq 32.70 Hz
        X"0017A7",  -- MIDI Note 25, Freq 34.65 Hz
        X"00190F",  -- MIDI Note 26, Freq 36.71 Hz
        X"001A8C",  -- MIDI Note 27, Freq 38.89 Hz
        X"001C20",  -- MIDI Note 28, Freq 41.20 Hz
        X"001DCD",  -- MIDI Note 29, Freq 43.65 Hz
        X"001F92",  -- MIDI Note 30, Freq 46.25 Hz
        X"002173",  -- MIDI Note 31, Freq 49.00 Hz
        X"002370",  -- MIDI Note 32, Freq 51.91 Hz
        X"00258B",  -- MIDI Note 33, Freq 55.00 Hz
        X"0027C7",  -- MIDI Note 34, Freq 58.27 Hz
        X"002A25",  -- MIDI Note 35, Freq 61.74 Hz
        X"002CA6",  -- MIDI Note 36, Freq 65.41 Hz
        X"002F4E",  -- MIDI Note 37, Freq 69.30 Hz
        X"00321E",  -- MIDI Note 38, Freq 73.42 Hz
        X"003519",  -- MIDI Note 39, Freq 77.78 Hz
        X"003841",  -- MIDI Note 40, Freq 82.41 Hz
        X"003B9A",  -- MIDI Note 41, Freq 87.31 Hz
        X"003F25",  -- MIDI Note 42, Freq 92.50 Hz
        X"0042E6",  -- MIDI Note 43, Freq 98.00 Hz
        X"0046E0",  -- MIDI Note 44, Freq 103.83 Hz
        X"004B17",  -- MIDI Note 45, Freq 110.00 Hz
        X"004F8F",  -- MIDI Note 46, Freq 116.54 Hz
        X"00544A",  -- MIDI Note 47, Freq 123.47 Hz
        X"00594D",  -- MIDI Note 48, Freq 130.81 Hz
        X"005E9C",  -- MIDI Note 49, Freq 138.59 Hz
        X"00643C",  -- MIDI Note 50, Freq 146.83 Hz
        X"006A32",  -- MIDI Note 51, Freq 155.56 Hz
        X"007083",  -- MIDI Note 52, Freq 164.81 Hz
        X"007734",  -- MIDI Note 53, Freq 174.61 Hz
        X"007E4A",  -- MIDI Note 54, Freq 185.00 Hz
        X"0085CD",  -- MIDI Note 55, Freq 196.00 Hz
        X"008DC1",  -- MIDI Note 56, Freq 207.65 Hz
        X"00962F",  -- MIDI Note 57, Freq 220.00 Hz
        X"009F1E",  -- MIDI Note 58, Freq 233.08 Hz
        X"00A894",  -- MIDI Note 59, Freq 246.94 Hz
        X"00B29A",  -- MIDI Note 60, Freq 261.63 Hz
        X"00BD39",  -- MIDI Note 61, Freq 277.18 Hz
        X"00C879",  -- MIDI Note 62, Freq 293.66 Hz
        X"00D465",  -- MIDI Note 63, Freq 311.13 Hz
        X"00E106",  -- MIDI Note 64, Freq 329.63 Hz
        X"00EE68",  -- MIDI Note 65, Freq 349.23 Hz
        X"00FC95",  -- MIDI Note 66, Freq 369.99 Hz
        X"010B9A",  -- MIDI Note 67, Freq 392.00 Hz
        X"011B83",  -- MIDI Note 68, Freq 415.30 Hz
        X"012C5F",  -- MIDI Note 69, Freq 440.00 Hz
        X"013E3C",  -- MIDI Note 70, Freq 466.16 Hz
        X"015128",  -- MIDI Note 71, Freq 493.88 Hz
        X"016534",  -- MIDI Note 72, Freq 523.25 Hz
        X"017A72",  -- MIDI Note 73, Freq 554.37 Hz
        X"0190F3",  -- MIDI Note 74, Freq 587.33 Hz
        X"01A8CA",  -- MIDI Note 75, Freq 622.25 Hz
        X"01C20D",  -- MIDI Note 76, Freq 659.26 Hz
        X"01DCD0",  -- MIDI Note 77, Freq 698.46 Hz
        X"01F92A",  -- MIDI Note 78, Freq 739.99 Hz
        X"021734",  -- MIDI Note 79, Freq 783.99 Hz
        X"023707",  -- MIDI Note 80, Freq 830.61 Hz
        X"0258BF",  -- MIDI Note 81, Freq 880.00 Hz
        X"027C78",  -- MIDI Note 82, Freq 932.33 Hz
        X"02A250",  -- MIDI Note 83, Freq 987.77 Hz
        X"02CA69",  -- MIDI Note 84, Freq 1046.50 Hz
        X"02F4E4",  -- MIDI Note 85, Freq 1108.73 Hz
        X"0321E6",  -- MIDI Note 86, Freq 1174.66 Hz
        X"035195",  -- MIDI Note 87, Freq 1244.51 Hz
        X"03841A",  -- MIDI Note 88, Freq 1318.51 Hz
        X"03B9A0",  -- MIDI Note 89, Freq 1396.91 Hz
        X"03F254",  -- MIDI Note 90, Freq 1479.98 Hz
        X"042E68",  -- MIDI Note 91, Freq 1567.98 Hz
        X"046E0F",  -- MIDI Note 92, Freq 1661.22 Hz
        X"04B17E",  -- MIDI Note 93, Freq 1760.00 Hz
        X"04F8F0",  -- MIDI Note 94, Freq 1864.66 Hz
        X"0544A1",  -- MIDI Note 95, Freq 1975.53 Hz
        X"0594D3",  -- MIDI Note 96, Freq 2093.00 Hz
        X"05E9C9",  -- MIDI Note 97, Freq 2217.46 Hz
        X"0643CD",  -- MIDI Note 98, Freq 2349.32 Hz
        X"06A32B",  -- MIDI Note 99, Freq 2489.02 Hz
        X"070834",  -- MIDI Note 100, Freq 2637.02 Hz
        X"077340",  -- MIDI Note 101, Freq 2793.83 Hz
        X"07E4A9",  -- MIDI Note 102, Freq 2959.96 Hz
        X"085CD1",  -- MIDI Note 103, Freq 3135.96 Hz
        X"08DC1E",  -- MIDI Note 104, Freq 3322.44 Hz
        X"0962FC",  -- MIDI Note 105, Freq 3520.00 Hz
        X"09F1E0",  -- MIDI Note 106, Freq 3729.31 Hz
        X"0A8942",  -- MIDI Note 107, Freq 3951.07 Hz
        X"0B29A6",  -- MIDI Note 108, Freq 4186.01 Hz
        X"0BD392",  -- MIDI Note 109, Freq 4434.92 Hz
        X"0C879A",  -- MIDI Note 110, Freq 4698.64 Hz
        X"0D4656",  -- MIDI Note 111, Freq 4978.03 Hz
        X"0E1069",  -- MIDI Note 112, Freq 5274.04 Hz
        X"0EE680",  -- MIDI Note 113, Freq 5587.65 Hz
        X"0FC953",  -- MIDI Note 114, Freq 5919.91 Hz
        X"10B9A2",  -- MIDI Note 115, Freq 6271.93 Hz
        X"11B83C",  -- MIDI Note 116, Freq 6644.88 Hz
        X"12C5F9",  -- MIDI Note 117, Freq 7040.00 Hz
        X"13E3C0",  -- MIDI Note 118, Freq 7458.62 Hz
        X"151285",  -- MIDI Note 119, Freq 7902.13 Hz
        X"16534C",  -- MIDI Note 120, Freq 8372.02 Hz
        X"17A725",  -- MIDI Note 121, Freq 8869.84 Hz
        X"190F34",  -- MIDI Note 122, Freq 9397.27 Hz
        X"1A8CAC",  -- MIDI Note 123, Freq 9956.06 Hz
        X"1C20D2",  -- MIDI Note 124, Freq 10548.08 Hz
        X"1DCD01",  -- MIDI Note 125, Freq 11175.30 Hz
        X"1F92A6",  -- MIDI Note 126, Freq 11839.82 Hz
        X"217345"  -- MIDI Note 127, Freq 12543.85 Hz
    );
end package body midi_lut_pkg;
